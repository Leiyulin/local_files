// this file is a *top file* of ctrl block
module mac_ctrl #
()
();

endmodule
