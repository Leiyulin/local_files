module phy_top#()
();

endmodule

PHY registers definition
32 registers
register 