module phy_top#()
();

endmodule